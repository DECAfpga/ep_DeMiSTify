../hdl/ctrl/demistify_config_pkg.vhd